`define IDX32(x) (((x)+1)*(32)-1):((x)*(32))
`define IDX8(x) (((x)+1)*(8)-1):((x)*(8))
`define BASE_VERSION 2
`define REVIS_ID 51
`define MF_PAR_ADD

module sha256_core(
	input i_clk,
	input i_rst_n,
	input [6:0] i_w_addr,
	input [7:0]	i_data8,
	input i_we,
	output o_irq,
	output reg [7:0] o_data_mux
);

	localparam START_W_MEM_ADDR = 0;
	localparam END_W_MEM_ADDR = 63;
	localparam WHO_AM_I = 7'd64;
	localparam STATUS_REG = 7'd65;
	localparam REVISION = 7'd66;
	localparam DAY = 7'd67;
	localparam MONTH = 7'd68;
	localparam YEAR = 7'd69;
	localparam WHO_AM_I_DATA = 7'd7;
	localparam REVISION_DATA = 8'd51;
	localparam DAY_DATA = 8'd19;
	localparam MONTH_DATA = 8'd03;
	localparam YEAR_DATA = 8'd19;
	localparam DIGEST_START_ADDR = 70;
	localparam DIGEST_END_ADDR = 101;

	`define ROUNDS4
	//`define ROUNDS16

	//16 addresses left empty
	localparam HASH_INIT = 256'h6a09e667_bb67ae85_3c6ef372_a54ff53a_510e527f_9b05688c_1f83d9ab_5be0cd19;

	// FSM states
    parameter   INIT = 2'd0,
                ROUND = 2'd1,
                MATH = 2'd2,
                OUT = 2'd3;

	reg [255:0] r_variables, r_variables_in; //a, b, c, d, e, f, g, h 
	reg [511:0] r_words; //W0, W1, W2 ... W15 in terms of FIPS
	reg [6:0] r_round, r_coef;
	reg [7:0] r_status; //r_status = {2'd0, r_state, completed, run, ready, start} // [7:1]read only [0] write accessable
	reg completed, run_signal, do_math;
	
	//variables indexing
	//wire [31:0] sum0_out, sum1_out, sigm0_out, sigm1_out, ch_out, maj_out, Kt_out;
	//wire [31:0] adder_wire_t1_1, adder_wire_t1_2, adder_wire_t1_3, t1, t2, adder_wire_word_1, adder_wire_word_2, new_word, new_a, new_e;
	wire [7:0] o_data_h;
	
	assign o_irq = completed;
	assign o_data_h = r_variables[(i_w_addr-DIGEST_START_ADDR) * 8 +: 8];

	// SPI data access
	always @* begin : data_access
		o_data_mux = 8'd0;
		if((i_w_addr >= 0) & (i_w_addr <= END_W_MEM_ADDR)) begin
			//o_data_mux = 8'd0;
		end else if (i_w_addr == WHO_AM_I) begin
			o_data_mux = WHO_AM_I_DATA;
		end else if (i_w_addr == STATUS_REG) begin
			o_data_mux = r_status;
		end else if(i_w_addr == REVISION) begin
			o_data_mux = REVISION_DATA;
		end else if(i_w_addr == DAY) begin
			o_data_mux = DAY_DATA;
		end else if(i_w_addr == MONTH) begin
			o_data_mux = MONTH_DATA;
		end else if(i_w_addr == YEAR) begin
			o_data_mux = YEAR_DATA;
		end else if ((i_w_addr >= DIGEST_START_ADDR) & (i_w_addr <= DIGEST_END_ADDR)) begin
			o_data_mux = o_data_h;
		end else if(i_w_addr > DIGEST_END_ADDR) begin
			o_data_mux = 8'haa;
		end
	end

    always @ (posedge i_clk or negedge i_rst_n) begin : hash_control_reg
        if(!i_rst_n) begin
            r_round <= 7'd0;
	    	r_coef <= 7'd0;
            r_status <= 8'd0;
			r_variables_in <= HASH_INIT;
        end else begin
        	if(i_we) begin
        		if(i_w_addr == STATUS_REG) begin
        			r_status <= i_data8[0];	
        		end
			end else begin
				case(r_status[5:4])
                	INIT: begin
                    	if(r_status[0]) begin
                        	r_status[5:4] <= ROUND;
                        	r_status[3:0] <= 4'b0100; //set start
							r_coef <= 7'd1;
							r_variables_in <= HASH_INIT;
                        end else begin
							r_coef <= 7'd0;
                        	r_status[3:0] <= 4'b0010; // ready
                        end
                	end
                	ROUND: begin
                		r_round <= r_round + 7'd8;
						r_coef <= r_coef + 7'd8;
						if(r_round == 7'd56) begin
                    		r_status[5:4] <= MATH;
                    		r_round <= 7'd0;
                    	end
                	end
                	MATH: begin
                		r_status[5:4] <= OUT;
                	end
                	OUT: begin
                		r_status <= 8'b0000_1010;
                		if(r_status[0]) begin
                			r_status[5:4] <= INIT;
                		end
                	end
                	default: begin end
            	endcase
			end             
        end
    end

    always @(*) begin : hash_control_comb
    	run_signal = 1'b0;
    	completed = 1'b0;
    	do_math = 1'b0;
    	case (r_status[5:4])
    		INIT: begin	end
    		ROUND: run_signal = 1'b1;
    		MATH: do_math = 1'b1;
    		OUT: completed = 1'b1;
    		default : /* default */;
    	endcase
    end

	// wire [255:0] variables_out_end;
	// wire [511:0] words_out_end;
	// wire [255:0] variables_out [0:ROUNDS-1];
	// wire [255:0] words_out [0:ROUNDS-1];

	// genvar i;
	// generate
	// 	for (i = 0; i < ROUNDS; i = i + 1) begin : HASHERS
	// 		if(i == 0) begin
	// 			sha256_digester_comb inst_sh (i_clk, r_round + i, r_variables, variables_out[i], r_words, words_out[i]);
	// 		end else if (i<ROUNDS-1) begin
	// 			sha256_digester_comb inst_sh (i_clk, r_round + i, variables_out[i-1], variables_out[i], words_out[i-1], words_out[i]);
	// 		end else begin
	// 			sha256_digester_comb inst_sh (i_clk, r_round + i, variables_out[i-1], variables_out_end, words_out[i-1], words_out_end);
	// 		end
	// 	end
	// endgenerate

	// Wires for round data transfer
	wire [255:0] variables_out1, variables_out2, variables_out3, variables_out4, variables_out5, variables_out6, variables_out7, variables_out8;
	wire [511:0] words_out1, words_out2, words_out3, words_out4, words_out5, words_out6, words_out7, words_out8;
	wire [255:0] variables_out9, variables_out10, variables_out11, variables_out12, variables_out13, variables_out14, variables_out15, variables_out16,variables_out_end;
	wire [511:0] words_out9, words_out10, words_out11, words_out12, words_out13, words_out14, words_out15, words_out16, words_out_end;
	wire [31:0] var_a, var_b, var_c, var_d, var_e, var_f, var_h, var_g;

	//Combinational cores
	
	sha256_digester_comb inst_sh1 (i_clk, r_round, 			 r_variables, variables_out1,    r_words, words_out1);
	sha256_digester_comb inst_sh2 (i_clk, r_round + 7'd1, variables_out1, variables_out2, words_out1, words_out2);
	sha256_digester_comb inst_sh3 (i_clk, r_round + 7'd2, variables_out2, variables_out3, words_out2, words_out3);
	sha256_digester_comb inst_sh4 (i_clk, r_round + 7'd3, variables_out3, variables_out4, words_out3, words_out4);

	`ifdef ROUNDS8
	sha256_digester_comb inst_sh5 (i_clk, r_round + 7'd4, variables_out4, variables_out5, words_out4, words_out5);
	sha256_digester_comb inst_sh6 (i_clk, r_round + 7'd5, variables_out5, variables_out6, words_out5, words_out6);
	sha256_digester_comb inst_sh7 (i_clk, r_round + 7'd6, variables_out6, variables_out7, words_out6, words_out7);
	sha256_digester_comb inst_sh8 (i_clk, r_round + 7'd7, variables_out7, variables_out8, words_out7, words_out8);
	`endif

	`ifdef ROUNDS16
	sha256_digester_comb inst_sh5 (i_clk, r_round + 7'd4, variables_out4, variables_out5, words_out4, words_out5);
	sha256_digester_comb inst_sh6 (i_clk, r_round + 7'd5, variables_out5, variables_out6, words_out5, words_out6);
	sha256_digester_comb inst_sh7 (i_clk, r_round + 7'd6, variables_out6, variables_out7, words_out6, words_out7);
	sha256_digester_comb inst_sh8 (i_clk, r_round + 7'd7, variables_out7, variables_out8, words_out7, words_out8);
	sha256_digester_comb inst_sh9 (i_clk, r_round + 7'd8, variables_out8, variables_out9, words_out8, words_out9);
	sha256_digester_comb inst_sh10 (i_clk, r_round + 7'd9, variables_out9, variables_out10, words_out9, words_out10);
	sha256_digester_comb inst_sh11 (i_clk, r_round + 7'd10, variables_out10, variables_out11, words_out10, words_out11);
	sha256_digester_comb inst_sh12 (i_clk, r_round + 7'd11, variables_out11, variables_out12, words_out11, words_out12);
	sha256_digester_comb inst_sh13 (i_clk, r_round + 7'd12, variables_out12, variables_out13, words_out12, words_out13);
	sha256_digester_comb inst_sh14 (i_clk, r_round + 7'd13, variables_out13, variables_out14, words_out13, words_out14);
	sha256_digester_comb inst_sh15 (i_clk, r_round + 7'd14, variables_out14, variables_out15, words_out14, words_out15);
	sha256_digester_comb inst_sh16 (i_clk, r_round + 7'd15, variables_out15, variables_out16, words_out15, words_out16);
	`endif

	`ifdef ROUNDS16
		assign variables_out_end = variables_out16;
		assign words_out_end = words_out16;
	`else 
		`ifdef ROUNDS8
			assign variables_out_end = variables_out8;
			assign words_out_end = words_out8;
		`else
			assign variables_out_end = variables_out4;
		assign words_out_end = words_out4;
		`endif
	`endif


	always @(posedge i_clk or negedge i_rst_n) begin : hash_math
		if(!i_rst_n) begin
			//r_variables_in <= HASH_INIT;
			r_words <= 512'd0;
			r_variables <= HASH_INIT;
		end else begin
			if (i_we & !run_signal) begin
				if ((i_w_addr >= START_W_MEM_ADDR) & (i_w_addr < (END_W_MEM_ADDR + 1))) begin
					r_words[(i_w_addr - START_W_MEM_ADDR) * 8 +: 8] <= i_data8;
				end
			end else if(run_signal & !i_we) begin : hash_computing
				r_words <= words_out_end;
				r_variables <= variables_out_end;
			end
			if(do_math) begin
				r_variables[`IDX32(7)] <= r_variables[`IDX32(7)] + r_variables_in[`IDX32(7)]; //<----------------- replace by adder module
				r_variables[`IDX32(6)] <= r_variables[`IDX32(6)] + r_variables_in[`IDX32(6)];	//replace by initial values for multiblock hash
				r_variables[`IDX32(5)] <= r_variables[`IDX32(5)] + r_variables_in[`IDX32(5)];
				r_variables[`IDX32(4)] <= r_variables[`IDX32(4)] + r_variables_in[`IDX32(4)];
				r_variables[`IDX32(3)] <= r_variables[`IDX32(3)] + r_variables_in[`IDX32(3)];
				r_variables[`IDX32(2)] <= r_variables[`IDX32(2)] + r_variables_in[`IDX32(2)];
				r_variables[`IDX32(1)] <= r_variables[`IDX32(1)] + r_variables_in[`IDX32(1)];
				r_variables[`IDX32(0)] <= r_variables[`IDX32(0)] + r_variables_in[`IDX32(0)];
			end
		end
	end
endmodule

module sha256_digester_comb (i_clk, r_coef, variables, o_variables, words, o_words);
	input i_clk;
	input [6:0] r_coef;
	input [511:0] words;
	input [255:0] variables;
	output [255:0] o_variables;
	output reg [511:0] o_words;

	wire [31:0] var_a = variables[`IDX32(7)];
	wire [31:0] var_b = variables[`IDX32(6)];
	wire [31:0] var_c = variables[`IDX32(5)];
	wire [31:0] var_d = variables[`IDX32(4)];
	wire [31:0] var_e = variables[`IDX32(3)];
	wire [31:0] var_f = variables[`IDX32(2)];
	wire [31:0] var_g = variables[`IDX32(1)];
	wire [31:0] var_h = variables[`IDX32(0)];
	reg [31:0] o_var_a, o_var_b, o_var_c, o_var_d, o_var_e, o_var_f, o_var_g, o_var_h;

	assign o_variables = {o_var_a, o_var_b, o_var_c, o_var_d, o_var_e, o_var_f, o_var_g, o_var_h};

	// SHA math and coef output
	wire [31:0] sum0_out, sum1_out, sigm0_out, sigm1_out, ch_out, maj_out, Kt_out;
	wire [31:0] new_word, new_a, new_e;
	//wire [31:0] adder_wire_t1_1, adder_wire_t1_2, adder_wire_t1_3, t1, t2, adder_wire_word_1, adder_wire_word_2, new_word, new_a, new_e;

	// `ifndef MF_PAR_ADD

	// //t1 adders, step 1
	// `ifdef ADD1
	// wire carryo1, carryo2, carryo3, carryo4, carryo5, carryo6, carryo7, carryo8, carryo9, carryo10;
	// wire [31:0] adder_wire_kt_ch, adder_wire_sum_wt, adder_wire_d_h, adder_wire_sum_wt_kt_ch, addw_maj_sum0, addw_sum_wt_kt_ch_h;
	// adder_32b_param st1_kt_ch (Kt_out, ch_out, 1'b0, carryo1, adder_wire_kt_ch);
	// adder_32b_param st1_sum_wt (sum1_out, words[`IDX32(15)], 1'b0, carryo2, adder_wire_sum_wt);
	// adder_32b_param st1_d_h (var_d, var_h, 1'b0, carryo3, adder_wire_d_h);

	// //t1 adders, step 2
	// adder_32b_param st2_sum_wt_kt_ch (adder_wire_kt_ch, adder_wire_sum_wt, 1'b0, carryo4, adder_wire_sum_wt_kt_ch);
	// adder_32b_param st2_all (adder_wire_sum_wt_kt_ch, adder_wire_d_h, 1'b0, carryo5, new_e);

	// //t1 adders, step 2 duplicate
	// adder_32b_param st2_a (adder_wire_sum_wt_kt_ch, var_h, 1'b0, carryo6, addw_sum_wt_kt_ch_h);
	// adder_32b_param st2_maj_sum0 (maj_out, sum0_out, 1'b0, carryo11, addw_maj_sum0);
	// adder_32b_param st2_a(addw_maj_sum0, addw_sum_wt_kt_ch_h, 1'b0, carryo12, new_a);

	// //new word adders
	// adder_32b_param inst_word_sigm1_rx_word (sigm1_out, words[`IDX32(6)], 1'b0, carryo8, adder_wire_word_1);
	// adder_32b_param inst_word_prev_sigm0 (adder_wire_word_1, sigm0_out, 1'b0, carryo9, adder_wire_word_2);
	// adder_32b_param inst_word_prev_words (adder_wire_word_2, words[`IDX32(15)], 1'b0, carryo10, new_word);
	// `endif

	// `ifdef ADD2
	// wire carryo1, carryo2, carryo3, carryo4, carryo5, carryo6, carryo7, carryo8, carryo9, carryo10;
	// wire [31:0] addw_kt_wt, adder_wire_sum_wt, adder_wire_d_h, adder_wire_sum_wt_kt_ch;

	// adder_32b_param add_kt_wt (Kt_out, words[`IDX32(15)], 1'b0, carryo1, addw_kt_wt);
	// adder_32b_param add_sum_ch (sum1_out, ch_out, 1'b0, carryo2, addw_sum_ch);
	// adder_32b_param add_d_h (var_d, var_h, 1'b0, carryo3, addw_d_h);

	// //t1 adders, step 2
	// adder_32b_param add_kt_wt_sum_ch (addw_kt_wt, addw_sum_ch, 1'b0, carryo4, addw_kt_wt_sum_ch);
	// adder_32b_param st2_all (addw_kt_wt_sum_ch, addw_d_h, 1'b0, carryo5, new_e);
	
	// //t1 adders, step 2 duplicate
	// adder_32b_param st2_a (adder_wire_sum_wt_kt_ch, var_h, 1'b0, carryo6, addw_sum_wt_kt_ch_h);
	// adder_32b_param st2_maj_sum0 (maj_out, sum0_out, 1'b0, carryo11, addw_maj_sum0);
	// adder_32b_param st2_a(addw_maj_sum0, addw_sum_wt_kt_ch_h, 1'b0, carryo12, new_a);

	// //new word adders
	// adder_32b_param inst_word_sigm1_rx_word (sigm1_out, words[`IDX32(6)], 1'b0, carryo8, adder_wire_word_1);
	// adder_32b_param inst_word_prev_sigm0 (adder_wire_word_1, sigm0_out, 1'b0, carryo9, adder_wire_word_2);
	// adder_32b_param inst_word_prev_words (adder_wire_word_2, words[`IDX32(15)], 1'b0, carryo10, new_word);
	// `endif

	// `else

	`ifdef MODEL_TECH
	assign new_e = Kt_out + ch_out + sum1_out + words[`IDX32(15)] + var_h + var_d;
	assign new_a = Kt_out + ch_out + sum1_out + words[`IDX32(15)] + var_h + maj_out + sum0_out;
	assign new_word = sigm1_out + words[`IDX32(6)] + sigm0_out + words[`IDX32(15)];
	`else
	par_add_6	par_add_6_inst (
								.data0x (Kt_out),
								.data1x (ch_out),
								.data2x (sum1_out),
								.data3x (words[`IDX32(15)]),
								.data4x (var_h),
								.data5x (var_d),
								.result (new_e)
								);

	par_add_7	par_add_7_inst (
								.data0x (Kt_out),
								.data1x (ch_out),
								.data2x (sum1_out),
								.data3x (words[`IDX32(15)]),
								.data4x (var_h),
								.data5x (maj_out),
								.data6x (sum0_out),
								.result (new_a)
								);

	par_add_4	par_add_4_inst (
								.data0x (sigm1_out),
								.data1x (words[`IDX32(6)]),
								.data2x (sigm0_out),
								.data3x (words[`IDX32(15)]),
								.result (new_word)
								);
	`endif
	

	sum0 inst_sum0(.x(var_a), .y(sum0_out));
	sum1 inst_sum1(.x(var_e), .y(sum1_out));
	sigm0 inst_sigm0(.x(words[`IDX32(14)]), .y(sigm0_out));
	sigm1 inst_sigm1(.x(words[`IDX32(1)]), .y(sigm1_out));
	ch inst_ch(.x(var_e), .y(var_f), .z(var_g), .o(ch_out));
	maj inst_maj(.x(var_a), .y(var_b), .z(var_c), .o(maj_out));
	sha256_coefs inst_coef(.i_coef_num(r_coef), .o_coef_value(Kt_out));

	//sha256_coefs_clk inst_coef_clk(.i_coef_num(r_coef), .i_clk(i_clk), .o_coef_value(Kt_out));

	always @* begin : hash_math
			o_words = {words[479:0], new_word};  //shift right replaced with shift left! <----------------- critical
			o_var_a = new_a; 		// new a from adder instance
			o_var_b = var_a;		// new b
			o_var_c = var_b;		// new c
			o_var_d = var_c;		// new d
			o_var_e = new_e;		// new e from adder instance, highest delay here
			o_var_f = var_e;		// new f
			o_var_g = var_f;		// new g
			o_var_h = var_g;		// new h
	end
endmodule